module alu_control (
    input instruction 
)

endmodule