// instruction_memory.v
`timescale 1ns/1ps
`include "params.vh"

module imem (
/* verilator lint_off UNUSEDSIGNAL */
input wire [63:0] pc, // reads from PC
input wire clk,
output reg [31:0] instruction // reads from memory the instruction 

);
  localparam MEMSIZE = 1024; // 1024 Instructions ~ 1024*4 = 4Kib
  localparam INSTRUCTION_N = 8;
  reg [31:0] i_mem[0:MEMSIZE-1];

initial begin 
    // Using assembly generated by my minimal rust assembler (https://github.com/1957-001B/ArmAsm)
    i_mem[0] = 32'hd2800088;  // "MOVZ X8, #0x4"
    i_mem[1] = 32'hd2800020;  // "MOVZ X0, #0x1"
    i_mem[2] = 32'h58000081;  // "LDR X1, =message"
    i_mem[3] = 32'hd28001a2;  // "MOVZ X2, #0xD"
    i_mem[4] = 32'hd2800028;
    i_mem[5] = 32'hd2800000;
    i_mem[6] = 32'hd4000001;
    i_mem[7] = 32'hE1000070;   // HLT #0 

    for (integer i = INSTRUCTION_N; i < MEMSIZE; i = i+1) begin
      i_mem[i] = 32'hd540643f; // NOP
    end

  end

  always @(posedge clk) begin
    instruction <= i_mem[pc[11:2]]; // right shifted twice to align with the 4 bit instuctions (i.e divide by 4)
  end

endmodule
