module registers(
  input clk;
  input [63:0] data_in,
  input [4:0] addr_write,
  input [9:5] addr_read,
 )




