
`ifndef INSTRUCTIONS_VH
`define INSTRUCTIONS_VH
DEFINE INSTRUCTION_N = 6;
instruction [0] = 32'h0x88;
instruction [1] = 32'h0x0;
instruction [2] = 32'h0x80;
instruction [3] = 32'h0xd2;
instruction [4] = 32'h0x20;
instruction [5] = 32'h0x0;
instruction [6] = 32'h0x80;
instruction [7] = 32'h0xd2;
instruction [8] = 32'h0xa2;
instruction [9] = 32'h0x1;
instruction [10] = 32'h0x80;
instruction [11] = 32'h0xd2;
instruction [12] = 32'h0x28;
instruction [13] = 32'h0x0;
instruction [14] = 32'h0x80;
instruction [15] = 32'h0xd2;
instruction [16] = 32'h0x0;
instruction [17] = 32'h0x0;
instruction [18] = 32'h0x80;
instruction [19] = 32'h0xd2;
instruction [20] = 32'h0x0;
instruction [21] = 32'h0x0;
instruction [22] = 32'h0x0;
instruction [23] = 32'h0x0;
endif
