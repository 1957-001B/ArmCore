module dmem (
    input [63:0] address,
    input [63:0] Write_d,
    output [63:0] Read_d
)
endmodule