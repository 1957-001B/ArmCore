`ifndef PARAMS_VH
`define PARAMS_VH
localparam CBZ_OP  = 8'b10110100;
localparam MOVZ_OP = 9'b110100101;
localparam CMP_OP  = 11'b11101011001;
localparam SUB_OP  = 9'b110100010;
localparam ADD_OP  = 9'b100100010;
localparam B_OP    = 6'b000101;
`endif